module systolic_multiplier #(parameter p_WORD_WIDTH = 4)(
	input wire i_CLK,
	input wire [p_WORD_WIDTH-1:0] i_MULTIPLIER,
	input wire i_MULTIPLICAND,
	output wire o_OUTPUT
);

wire [p_WORD_WIDTH-1:0] w_CARRY_FEEDBACK;
wire [p_WORD_WIDTH-2:0] w_CELL_INTERCONNECT_RESULT;
wire [p_WORD_WIDTH-2:0] w_CELL_INTERCONNECT_BROADCAST;
systolic_mult_cell s0 (
	.i_CLK(i_CLK),
	.i_INPUT(i_MULTIPLICAND),
	.i_CARRY_IN(w_CARRY_FEEDBACK[0]),
	.i_WEIGHT(i_MULTIPLIER[0]),
	.i_ADJ_RESULT(w_CELL_INTERCONNECT_RESULT[0]),
	.o_INPUT_BROADCAST(w_CELL_INTERCONNECT_BROADCAST[0]),
	.o_CARRY_OUT(w_CARRY_FEEDBACK[0]),
	.o_OUTPUT(o_OUTPUT)
);
systolic_mult_cell s1 (
	.i_CLK(i_CLK),
	.i_INPUT(w_CELL_INTERCONNECT_BROADCAST[0]),
	.i_CARRY_IN(w_CARRY_FEEDBACK[1]),
	.i_WEIGHT(i_MULTIPLIER[1]),
	.i_ADJ_RESULT(w_CELL_INTERCONNECT_RESULT[1]),
	.o_INPUT_BROADCAST(w_CELL_INTERCONNECT_BROADCAST[1]),
	.o_CARRY_OUT(w_CARRY_FEEDBACK[1]),
	.o_OUTPUT(w_CELL_INTERCONNECT_RESULT[0])
);
systolic_mult_cell s2 (
	.i_CLK(i_CLK),
	.i_INPUT(w_CELL_INTERCONNECT_BROADCAST[1]),
	.i_CARRY_IN(w_CARRY_FEEDBACK[2]),
	.i_WEIGHT(i_MULTIPLIER[2]),
	.i_ADJ_RESULT(w_CELL_INTERCONNECT_RESULT[2]),
	.o_INPUT_BROADCAST(w_CELL_INTERCONNECT_BROADCAST[2]),
	.o_CARRY_OUT(w_CARRY_FEEDBACK[2]),
	.o_OUTPUT(w_CELL_INTERCONNECT_RESULT[1])
);
systolic_mult_cell s3 (
	.i_CLK(i_CLK),
	.i_INPUT(w_CELL_INTERCONNECT_BROADCAST[2]),
	.i_CARRY_IN(w_CARRY_FEEDBACK[3]),
	.i_WEIGHT(i_MULTIPLIER[3]),
	.i_ADJ_RESULT(),
	.o_INPUT_BROADCAST(),
	.o_CARRY_OUT(w_CARRY_FEEDBACK[3]),
	.o_OUTPUT(w_CELL_INTERCONNECT_RESULT[2])
);
endmodule
