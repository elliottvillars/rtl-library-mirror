
module simple_axi_slave(
);
//TODO: Add singals
endmodule
