module single_port_bram (
	input wire i_CLK,
	input wire i_WRITE_ENABLE,
	input wire i_READ_ENABLE,
	input wire i_ADDRESS,
	input wire i_WRITE_DATA,
	output reg o_READ_DATA
);
endmodule
