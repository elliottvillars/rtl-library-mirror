`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/09/2018 12:15:35 PM
// Design Name: 
// Module Name: HZ_Counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`default_nettype none
module static_clock_divider(
	input wire i_CLK,
	input wire i_RESET,
	input wire i_ENABLE,
	output reg o_ENABLE_OUT
);

parameter p_DIV_VALUE = 3;
reg [31:0] r_Count;
always @ (posedge(i_CLK)) //Counter
begin
	if (i_RESET == 1'b1)
	begin
		r_Count <= 32'b0;
	end
	else
	begin
		if(i_ENABLE == 1'b1) 
		begin
			if (r_Count >= p_DIV_VALUE)
				r_Count <= 32'b0;
			else
				r_Count <= r_Count + 1;
		end
		else
		begin
			r_Count <= 32'd0;
		end
	end
end

always @ (posedge(i_CLK)) //FF with comparator
begin
	if (i_RESET == 1'b1)
	begin
		o_ENABLE_OUT <= 1'b0;
	end
	else 
	begin
		if (r_Count == p_DIV_VALUE && i_ENABLE == 1) // if r_Count = 49999999 flip output
		begin
			o_ENABLE_OUT <= 1'b1;
		end
		else
		begin
			o_ENABLE_OUT <= 1'b0;
		end
	end
end

//TODO:Perform QA pass and reverify this module.
`ifdef FORMAL
	reg r_PAST_VALID;
	initial begin
		assume(r_Count == 0);
		assume(i_CLK == 0);
		assume(i_RESET == 1);
	end

	always@(posedge i_CLK)
	begin
		r_PAST_VALID = 1;
		assume(i_CLK != $past(i_CLK));
		if(r_PAST_VALID == 1 && $rose(i_CLK))
		begin
			if($past(i_RESET) == 1)
			begin
				assert(r_Count == 0);
				assert(o_ENABLE_OUT == 0);
			end
			else
			begin
				if($stable(i_RESET) && $past(i_RESET) == 0)
				begin
					if($stable(i_ENABLE) && $past(i_ENABLE) == 1)
					begin
						if($past(r_Count) != p_DIV_VALUE)
							assert(o_ENABLE_OUT == 0);
						else
						begin
							assert(o_ENABLE_OUT == 1);
							assert(r_Count == 0);
						end
					end
				end
			end
		end
	end
`endif
endmodule
