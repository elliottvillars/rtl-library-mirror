module foo (
);
endmodule
