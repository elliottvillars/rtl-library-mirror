module foo (
	input i_CLK
);
`ifdef FORMAL
`endif
endmodule
